module top_module(
   zero
);// Module body starts after semicolon
	output zero;
endmodule
