module top_module( 
    input a, 
    input b, 
    output out );

    assign out = !(a^b);
    //Or
    //assign out = (((!a)&&(!b))||(a&&b));

endmodule
